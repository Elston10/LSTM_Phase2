// Corrected Tanh LUT for S7.8 Fixed-Point Format
// Input range: [0.25, 3.0] with step size 0.01
// Contains actual tanh(x) values, not linear progression

module tanh_lut_ram #(
    parameter WIDTH = 16,
    parameter ADDR_WIDTH = 9,
    parameter LUT_SIZE = 276
) (
    input  [ADDR_WIDTH-1:0] addr,
    output [WIDTH-1:0] tanh_out
);

    // LUT data array
    reg [WIDTH-1:0] tanh_lut [0:LUT_SIZE-1];
 initial begin   
    // Initialize LUT with ACTUAL tanh values
     tanh_lut[  0] = 16'h003F; // tanh(0.25)
    tanh_lut[  1] = 16'h0041; // tanh(0.26)
    tanh_lut[  2] = 16'h0043; // tanh(0.27)
    tanh_lut[  3] = 16'h0046; // tanh(0.28)
    tanh_lut[  4] = 16'h0048; // tanh(0.29)
    tanh_lut[  5] = 16'h004B; // tanh(0.30)
    tanh_lut[  6] = 16'h004D; // tanh(0.31)
    tanh_lut[  7] = 16'h004F; // tanh(0.32)
    tanh_lut[  8] = 16'h0052; // tanh(0.33)
    tanh_lut[  9] = 16'h0054; // tanh(0.34)
    tanh_lut[ 10] = 16'h0056; // tanh(0.35)
    tanh_lut[ 11] = 16'h0058; // tanh(0.36)
    tanh_lut[ 12] = 16'h005B; // tanh(0.37)
    tanh_lut[ 13] = 16'h005D; // tanh(0.38)
    tanh_lut[ 14] = 16'h005F; // tanh(0.39)
    tanh_lut[ 15] = 16'h0061; // tanh(0.40)
    tanh_lut[ 16] = 16'h0063; // tanh(0.41)
    tanh_lut[ 17] = 16'h0066; // tanh(0.42)
    tanh_lut[ 18] = 16'h0068; // tanh(0.43)
    tanh_lut[ 19] = 16'h006A; // tanh(0.44)
    tanh_lut[ 20] = 16'h006C; // tanh(0.45)
    tanh_lut[ 21] = 16'h006E; // tanh(0.46)
    tanh_lut[ 22] = 16'h0070; // tanh(0.47)
    tanh_lut[ 23] = 16'h0072; // tanh(0.48)
    tanh_lut[ 24] = 16'h0074; // tanh(0.49)
    tanh_lut[ 25] = 16'h0076; // tanh(0.50)
    tanh_lut[ 26] = 16'h0078; // tanh(0.51)
    tanh_lut[ 27] = 16'h007A; // tanh(0.52)
    tanh_lut[ 28] = 16'h007C; // tanh(0.53)
    tanh_lut[ 29] = 16'h007E; // tanh(0.54)
    tanh_lut[ 30] = 16'h0080; // tanh(0.55)
    tanh_lut[ 31] = 16'h0082; // tanh(0.56)
    tanh_lut[ 32] = 16'h0084; // tanh(0.57)
    tanh_lut[ 33] = 16'h0086; // tanh(0.58)
    tanh_lut[ 34] = 16'h0088; // tanh(0.59)
    tanh_lut[ 35] = 16'h0089; // tanh(0.60)
    tanh_lut[ 36] = 16'h008B; // tanh(0.61)
    tanh_lut[ 37] = 16'h008D; // tanh(0.62)
    tanh_lut[ 38] = 16'h008F; // tanh(0.63)
    tanh_lut[ 39] = 16'h0091; // tanh(0.64)
    tanh_lut[ 40] = 16'h0092; // tanh(0.65)
    tanh_lut[ 41] = 16'h0094; // tanh(0.66)
    tanh_lut[ 42] = 16'h0096; // tanh(0.67)
    tanh_lut[ 43] = 16'h0097; // tanh(0.68)
    tanh_lut[ 44] = 16'h0099; // tanh(0.69)
    tanh_lut[ 45] = 16'h009B; // tanh(0.70)
    tanh_lut[ 46] = 16'h009C; // tanh(0.71)
    tanh_lut[ 47] = 16'h009E; // tanh(0.72)
    tanh_lut[ 48] = 16'h00A0; // tanh(0.73)
    tanh_lut[ 49] = 16'h00A1; // tanh(0.74)
    tanh_lut[ 50] = 16'h00A3; // tanh(0.75)
    tanh_lut[ 51] = 16'h00A4; // tanh(0.76)
    tanh_lut[ 52] = 16'h00A6; // tanh(0.77)
    tanh_lut[ 53] = 16'h00A7; // tanh(0.78)
    tanh_lut[ 54] = 16'h00A9; // tanh(0.79)
    tanh_lut[ 55] = 16'h00AA; // tanh(0.80)
    tanh_lut[ 56] = 16'h00AB; // tanh(0.81)
    tanh_lut[ 57] = 16'h00AD; // tanh(0.82)
    tanh_lut[ 58] = 16'h00AE; // tanh(0.83)
    tanh_lut[ 59] = 16'h00B0; // tanh(0.84)
    tanh_lut[ 60] = 16'h00B1; // tanh(0.85)
    tanh_lut[ 61] = 16'h00B2; // tanh(0.86)
    tanh_lut[ 62] = 16'h00B4; // tanh(0.87)
    tanh_lut[ 63] = 16'h00B5; // tanh(0.88)
    tanh_lut[ 64] = 16'h00B6; // tanh(0.89)
    tanh_lut[ 65] = 16'h00B7; // tanh(0.90)
    tanh_lut[ 66] = 16'h00B9; // tanh(0.91)
    tanh_lut[ 67] = 16'h00BA; // tanh(0.92)
    tanh_lut[ 68] = 16'h00BB; // tanh(0.93)
    tanh_lut[ 69] = 16'h00BC; // tanh(0.94)
    tanh_lut[ 70] = 16'h00BD; // tanh(0.95)
    tanh_lut[ 71] = 16'h00BF; // tanh(0.96)
    tanh_lut[ 72] = 16'h00C0; // tanh(0.97)
    tanh_lut[ 73] = 16'h00C1; // tanh(0.98)
    tanh_lut[ 74] = 16'h00C2; // tanh(0.99)
    tanh_lut[ 75] = 16'h00C3; // tanh(1.00)
    tanh_lut[ 76] = 16'h00C4; // tanh(1.01)
    tanh_lut[ 77] = 16'h00C5; // tanh(1.02)
    tanh_lut[ 78] = 16'h00C6; // tanh(1.03)
    tanh_lut[ 79] = 16'h00C7; // tanh(1.04)
    tanh_lut[ 80] = 16'h00C8; // tanh(1.05)
    tanh_lut[ 81] = 16'h00C9; // tanh(1.06)
    tanh_lut[ 82] = 16'h00CA; // tanh(1.07)
    tanh_lut[ 83] = 16'h00CB; // tanh(1.08)
    tanh_lut[ 84] = 16'h00CC; // tanh(1.09)
    tanh_lut[ 85] = 16'h00CD; // tanh(1.10)
    tanh_lut[ 86] = 16'h00CE; // tanh(1.11)
    tanh_lut[ 87] = 16'h00CF; // tanh(1.12)
    tanh_lut[ 88] = 16'h00D0; // tanh(1.13)
    tanh_lut[ 89] = 16'h00D0; // tanh(1.14)
    tanh_lut[ 90] = 16'h00D1; // tanh(1.15)
    tanh_lut[ 91] = 16'h00D2; // tanh(1.16)
    tanh_lut[ 92] = 16'h00D3; // tanh(1.17)
    tanh_lut[ 93] = 16'h00D4; // tanh(1.18)
    tanh_lut[ 94] = 16'h00D5; // tanh(1.19)
    tanh_lut[ 95] = 16'h00D5; // tanh(1.20)
    tanh_lut[ 96] = 16'h00D6; // tanh(1.21)
    tanh_lut[ 97] = 16'h00D7; // tanh(1.22)
    tanh_lut[ 98] = 16'h00D8; // tanh(1.23)
    tanh_lut[ 99] = 16'h00D8; // tanh(1.24)
    tanh_lut[100] = 16'h00D9; // tanh(1.25)
    tanh_lut[101] = 16'h00DA; // tanh(1.26)
    tanh_lut[102] = 16'h00DB; // tanh(1.27)
    tanh_lut[103] = 16'h00DB; // tanh(1.28)
    tanh_lut[104] = 16'h00DC; // tanh(1.29)
    tanh_lut[105] = 16'h00DD; // tanh(1.30)
    tanh_lut[106] = 16'h00DD; // tanh(1.31)
    tanh_lut[107] = 16'h00DE; // tanh(1.32)
    tanh_lut[108] = 16'h00DF; // tanh(1.33)
    tanh_lut[109] = 16'h00DF; // tanh(1.34)
    tanh_lut[110] = 16'h00E0; // tanh(1.35)
    tanh_lut[111] = 16'h00E0; // tanh(1.36)
    tanh_lut[112] = 16'h00E1; // tanh(1.37)
    tanh_lut[113] = 16'h00E2; // tanh(1.38)
    tanh_lut[114] = 16'h00E2; // tanh(1.39)
    tanh_lut[115] = 16'h00E3; // tanh(1.40)
    tanh_lut[116] = 16'h00E3; // tanh(1.41)
    tanh_lut[117] = 16'h00E4; // tanh(1.42)
    tanh_lut[118] = 16'h00E4; // tanh(1.43)
    tanh_lut[119] = 16'h00E5; // tanh(1.44)
    tanh_lut[120] = 16'h00E5; // tanh(1.45)
    tanh_lut[121] = 16'h00E6; // tanh(1.46)
    tanh_lut[122] = 16'h00E6; // tanh(1.47)
    tanh_lut[123] = 16'h00E7; // tanh(1.48)
    tanh_lut[124] = 16'h00E7; // tanh(1.49)
    tanh_lut[125] = 16'h00E8; // tanh(1.50)
    tanh_lut[126] = 16'h00E8; // tanh(1.51)
    tanh_lut[127] = 16'h00E9; // tanh(1.52)
    tanh_lut[128] = 16'h00E9; // tanh(1.53)
    tanh_lut[129] = 16'h00EA; // tanh(1.54)
    tanh_lut[130] = 16'h00EA; // tanh(1.55)
    tanh_lut[131] = 16'h00EA; // tanh(1.56)
    tanh_lut[132] = 16'h00EB; // tanh(1.57)
    tanh_lut[133] = 16'h00EB; // tanh(1.58)
    tanh_lut[134] = 16'h00EC; // tanh(1.59)
    tanh_lut[135] = 16'h00EC; // tanh(1.60)
    tanh_lut[136] = 16'h00EC; // tanh(1.61)
    tanh_lut[137] = 16'h00ED; // tanh(1.62)
    tanh_lut[138] = 16'h00ED; // tanh(1.63)
    tanh_lut[139] = 16'h00ED; // tanh(1.64)
    tanh_lut[140] = 16'h00EE; // tanh(1.65)
    tanh_lut[141] = 16'h00EE; // tanh(1.66)
    tanh_lut[142] = 16'h00EE; // tanh(1.67)
    tanh_lut[143] = 16'h00EF; // tanh(1.68)
    tanh_lut[144] = 16'h00EF; // tanh(1.69)
    tanh_lut[145] = 16'h00EF; // tanh(1.70)
    tanh_lut[146] = 16'h00F0; // tanh(1.71)
    tanh_lut[147] = 16'h00F0; // tanh(1.72)
    tanh_lut[148] = 16'h00F0; // tanh(1.73)
    tanh_lut[149] = 16'h00F1; // tanh(1.74)
    tanh_lut[150] = 16'h00F1; // tanh(1.75)
    tanh_lut[151] = 16'h00F1; // tanh(1.76)
    tanh_lut[152] = 16'h00F2; // tanh(1.77)
    tanh_lut[153] = 16'h00F2; // tanh(1.78)
    tanh_lut[154] = 16'h00F2; // tanh(1.79)
    tanh_lut[155] = 16'h00F2; // tanh(1.80)
    tanh_lut[156] = 16'h00F3; // tanh(1.81)
    tanh_lut[157] = 16'h00F3; // tanh(1.82)
    tanh_lut[158] = 16'h00F3; // tanh(1.83)
    tanh_lut[159] = 16'h00F3; // tanh(1.84)
    tanh_lut[160] = 16'h00F4; // tanh(1.85)
    tanh_lut[161] = 16'h00F4; // tanh(1.86)
    tanh_lut[162] = 16'h00F4; // tanh(1.87)
    tanh_lut[163] = 16'h00F4; // tanh(1.88)
    tanh_lut[164] = 16'h00F5; // tanh(1.89)
    tanh_lut[165] = 16'h00F5; // tanh(1.90)
    tanh_lut[166] = 16'h00F5; // tanh(1.91)
    tanh_lut[167] = 16'h00F5; // tanh(1.92)
    tanh_lut[168] = 16'h00F5; // tanh(1.93)
    tanh_lut[169] = 16'h00F6; // tanh(1.94)
    tanh_lut[170] = 16'h00F6; // tanh(1.95)
    tanh_lut[171] = 16'h00F6; // tanh(1.96)
    tanh_lut[172] = 16'h00F6; // tanh(1.97)
    tanh_lut[173] = 16'h00F6; // tanh(1.98)
    tanh_lut[174] = 16'h00F7; // tanh(1.99)
    tanh_lut[175] = 16'h00F7; // tanh(2.00)
    tanh_lut[176] = 16'h00F7; // tanh(2.01)
    tanh_lut[177] = 16'h00F7; // tanh(2.02)
    tanh_lut[178] = 16'h00F7; // tanh(2.03)
    tanh_lut[179] = 16'h00F7; // tanh(2.04)
    tanh_lut[180] = 16'h00F8; // tanh(2.05)
    tanh_lut[181] = 16'h00F8; // tanh(2.06)
    tanh_lut[182] = 16'h00F8; // tanh(2.07)
    tanh_lut[183] = 16'h00F8; // tanh(2.08)
    tanh_lut[184] = 16'h00F8; // tanh(2.09)
    tanh_lut[185] = 16'h00F8; // tanh(2.10)
    tanh_lut[186] = 16'h00F9; // tanh(2.11)
    tanh_lut[187] = 16'h00F9; // tanh(2.12)
    tanh_lut[188] = 16'h00F9; // tanh(2.13)
    tanh_lut[189] = 16'h00F9; // tanh(2.14)
    tanh_lut[190] = 16'h00F9; // tanh(2.15)
    tanh_lut[191] = 16'h00F9; // tanh(2.16)
    tanh_lut[192] = 16'h00F9; // tanh(2.17)
    tanh_lut[193] = 16'h00FA; // tanh(2.18)
    tanh_lut[194] = 16'h00FA; // tanh(2.19)
    tanh_lut[195] = 16'h00FA; // tanh(2.20)
    tanh_lut[196] = 16'h00FA; // tanh(2.21)
    tanh_lut[197] = 16'h00FA; // tanh(2.22)
    tanh_lut[198] = 16'h00FA; // tanh(2.23)
    tanh_lut[199] = 16'h00FA; // tanh(2.24)
    tanh_lut[200] = 16'h00FA; // tanh(2.25)
    tanh_lut[201] = 16'h00FA; // tanh(2.26)
    tanh_lut[202] = 16'h00FB; // tanh(2.27)
    tanh_lut[203] = 16'h00FB; // tanh(2.28)
    tanh_lut[204] = 16'h00FB; // tanh(2.29)
    tanh_lut[205] = 16'h00FB; // tanh(2.30)
    tanh_lut[206] = 16'h00FB; // tanh(2.31)
    tanh_lut[207] = 16'h00FB; // tanh(2.32)
    tanh_lut[208] = 16'h00FB; // tanh(2.33)
    tanh_lut[209] = 16'h00FB; // tanh(2.34)
    tanh_lut[210] = 16'h00FB; // tanh(2.35)
    tanh_lut[211] = 16'h00FB; // tanh(2.36)
    tanh_lut[212] = 16'h00FC; // tanh(2.37)
    tanh_lut[213] = 16'h00FC; // tanh(2.38)
    tanh_lut[214] = 16'h00FC; // tanh(2.39)
    tanh_lut[215] = 16'h00FC; // tanh(2.40)
    tanh_lut[216] = 16'h00FC; // tanh(2.41)
    tanh_lut[217] = 16'h00FC; // tanh(2.42)
    tanh_lut[218] = 16'h00FC; // tanh(2.43)
    tanh_lut[219] = 16'h00FC; // tanh(2.44)
    tanh_lut[220] = 16'h00FC; // tanh(2.45)
    tanh_lut[221] = 16'h00FC; // tanh(2.46)
    tanh_lut[222] = 16'h00FC; // tanh(2.47)
    tanh_lut[223] = 16'h00FC; // tanh(2.48)
    tanh_lut[224] = 16'h00FD; // tanh(2.49)
    tanh_lut[225] = 16'h00FD; // tanh(2.50)
    tanh_lut[226] = 16'h00FD; // tanh(2.51)
    tanh_lut[227] = 16'h00FD; // tanh(2.52)
    tanh_lut[228] = 16'h00FD; // tanh(2.53)
    tanh_lut[229] = 16'h00FD; // tanh(2.54)
    tanh_lut[230] = 16'h00FD; // tanh(2.55)
    tanh_lut[231] = 16'h00FD; // tanh(2.56)
    tanh_lut[232] = 16'h00FD; // tanh(2.57)
    tanh_lut[233] = 16'h00FD; // tanh(2.58)
    tanh_lut[234] = 16'h00FD; // tanh(2.59)
    tanh_lut[235] = 16'h00FD; // tanh(2.60)
    tanh_lut[236] = 16'h00FD; // tanh(2.61)
    tanh_lut[237] = 16'h00FD; // tanh(2.62)
    tanh_lut[238] = 16'h00FD; // tanh(2.63)
    tanh_lut[239] = 16'h00FD; // tanh(2.64)
    tanh_lut[240] = 16'h00FD; // tanh(2.65)
    tanh_lut[241] = 16'h00FE; // tanh(2.66)
    tanh_lut[242] = 16'h00FE; // tanh(2.67)
    tanh_lut[243] = 16'h00FE; // tanh(2.68)
    tanh_lut[244] = 16'h00FE; // tanh(2.69)
    tanh_lut[245] = 16'h00FE; // tanh(2.70)
    tanh_lut[246] = 16'h00FE; // tanh(2.71)
    tanh_lut[247] = 16'h00FE; // tanh(2.72)
    tanh_lut[248] = 16'h00FE; // tanh(2.73)
    tanh_lut[249] = 16'h00FE; // tanh(2.74)
    tanh_lut[250] = 16'h00FE; // tanh(2.75)
    tanh_lut[251] = 16'h00FE; // tanh(2.76)
    tanh_lut[252] = 16'h00FE; // tanh(2.77)
    tanh_lut[253] = 16'h00FE; // tanh(2.78)
    tanh_lut[254] = 16'h00FE; // tanh(2.79)
    tanh_lut[255] = 16'h00FE; // tanh(2.80)
    tanh_lut[256] = 16'h00FE; // tanh(2.81)
    tanh_lut[257] = 16'h00FE; // tanh(2.82)
    tanh_lut[258] = 16'h00FE; // tanh(2.83)
    tanh_lut[259] = 16'h00FE; // tanh(2.84)
    tanh_lut[260] = 16'h00FE; // tanh(2.85)
    tanh_lut[261] = 16'h00FE; // tanh(2.86)
    tanh_lut[262] = 16'h00FE; // tanh(2.87)
    tanh_lut[263] = 16'h00FE; // tanh(2.88)
    tanh_lut[264] = 16'h00FE; // tanh(2.89)
    tanh_lut[265] = 16'h00FE; // tanh(2.90)
    tanh_lut[266] = 16'h00FE; // tanh(2.91)
    tanh_lut[267] = 16'h00FF; // tanh(2.92)
    tanh_lut[268] = 16'h00FF; // tanh(2.93)
    tanh_lut[269] = 16'h00FF; // tanh(2.94)
    tanh_lut[270] = 16'h00FF; // tanh(2.95)
    tanh_lut[271] = 16'h00FF; // tanh(2.96)
    tanh_lut[272] = 16'h00FF; // tanh(2.97)
    tanh_lut[273] = 16'h00FF; // tanh(2.98)
    tanh_lut[274] = 16'h00FF; // tanh(2.99)
    tanh_lut[275] = 16'h00FF; // tanh(3.00)
end
    
    // Output assignment with bounds checking
    assign tanh_out = (addr < LUT_SIZE) ? tanh_lut[addr] : tanh_lut[LUT_SIZE-1];

endmodule